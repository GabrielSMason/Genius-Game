module reg_fpga
(
	clk_i,
	r_i,
	e_i,
	data_i,
	q_o,
	q3_o
);

localparam N = 64;
localparam N1 = 4;

input wire clk_i,r_i,e_i;
input wire [N-1:0]data_i;
output reg [N-1:0]q_o;
output reg [N1-1:0]q3_o;

always@(posedge clk_i or posedge r_i) begin 
	if(r_i) begin
		q_o <= 64'b0;
		q3_o <= 4'b0;
	end 
	else if (e_i) begin
		q_o <= data_i;
		q3_o <= data_i[63:60];
	end
end 

endmodule
