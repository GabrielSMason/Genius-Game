module decSeq00
(
	address_i,
	output_o
);

input [3:0]address_i;
output reg [3:0]output_o;

endmodule
